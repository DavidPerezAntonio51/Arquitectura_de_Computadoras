library ieee;
use ieee.std_logic_1164.all;

entity contring00 is port(
	
);
end entity;

architecture contring0 of contring00 is
begin

end architecture;