library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity barrelrotationLR is port(
	clks: in std_logic;
	ens: in std_logic;
	ins: in std_logic_vector(7 downto 0);
	outs: out std_logic_vector(7 downto 0);
	control: in std_logic_vector(3 downto 0)
);
end entity;

architecture barrelrotationLR0 of barrelrotationLR is
	signal srotation: std_logic_vector(7 downto 0);
	signal scontrol: std_logic_vector(3 downto 0);
begin
	pshift: process(clks)
	begin
	if(clks'event and clks = '1') then
		case ens is
			when '0' =>
				outs <= "00000000";
				srotation <= ins;
				scontrol<= "0000";
			when '1'=>
			if(scontrol<control)then
				scontrol <= scontrol + '1';
				-----------------
				srotation(7) <= srotation(0);
				srotation(6 downto 0) <= srotation(7 downto 1);
				outs <= srotation;
			else
				scontrol<=scontrol;
			end if;
			when others => null;
		end case;
	end if;
	end process pshift;
end architecture;